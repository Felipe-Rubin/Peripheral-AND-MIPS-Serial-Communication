-- PT_BR
------------------------------------------------------------------------
-- Autores : Felipe Rubin & Ariel Ril & Ney Calazans & Fernando Moraes
--
-- Email: felipe.rubin@acad.pucrs.br & ariel.ril@acad.pucrs.br & ney.calazans@pucrs.br & fernando.moraes@pucrs.br
--
-- T1 Organizacao e Arquitetura de Computadores II PUCRS 2017/2
--
-- Arquivo : System_tb.vhd
--
-- Descricao: Este arquivo representa o testbench do sistema. Este arquivo
-- foi gerado a partir de dois testbenches e hardware's implementados pelos professores
-- Ney Calazans e Fernando Moraes. Um testbench era da interface serial, enquanto outro
-- era o do MIPS. O trabalho em cima dele foi de criar um periferico
-- no testbench e um componente de hardware de logica de cola, assim montando
-- um sistema de transmissao e recepcao de dados.
------------------------------------------------------------------------
-- EN_US
------------------------------------------------------------------------
-- Authors : Felipe Rubin & Ariel Ril & Ney Calazans
--
-- Email: felipe.rubin@acad.pucrs.br & ariel.ril@acad.pucrs.br & ney.calazans@pucrs.br & fernando.moraes@pucrs.br
--
-- Assignment 1 Computer Organization and Design II PUCRS 2017/2
--
-- File : System_tb.vhd
--
-- Description: This file represents the system testbench. This file
-- was generated by two other testbenches and hardwares which were implemented by
-- professor Ney Calazans and professor Fernando Mores. One testebench was
--  for the serial interface, while the other was from MIPS. The assignment was 
-- to create a peripheral in the testbench and a hardware component of glue logic,
-- in order to create a system of transmission and reception of data.
------------------------------------------------------------------------


-------------------------------------------------------------------------
--
-- 32 bits PROCESSOR TESTBENCH    LITTLE  ENDIAN      13/october/2004
--
-- It must be observed that the processor is hold in reset
-- (reset <= '1') at the start of simulation, being activated
-- (reset <= '0') just after the end of the object file reading be the
-- testbench.
--
-- This testbench employs two memories, implying a HARVARD organization
--
-- Changes:
--	16/05/2012 (Ney Calazans)
--		- Corrected bug in memory filling during reset. The instruction
--		memory fill process, makes the processor produce "ce" signals to 
--		memory which ended up by filling data memory with rubbish at
--		the same time. To solve this, the first line of the data memory
--		Dce control signal generation was changed from 
--			--	ce='1' or go_d='1'	 to 
--			-- (ce='1' and reset/='1') or go_d='1'
--		- Also, there was a problem with the data memory write operation in
--		monocycle MIPS implementations: when multiple SW instructions
--		were issued one after the other, the write operation was executed
--		in two sets of memory positions at once after the first SW. To
--		solve this the data signal was removed from the memory write
--		process sensitivity list.
--	10/10/2015 (Ney Calazans)
--		- Signal bw from memory set to '1', since the CPU
--		does not generate it anymore.
--	28/10/2016 (Ney Calazans)
--		- Also, regX defs were changed to wiresX, to improve
--		code readability.
--	02/06/2017 (Ney Calazans) - bugfix
--		- tmp_address changed to int_address in the memory definition
--		-IN the definition of the memory read/write processes,
--		  CONV_INTEGER(low_address+3)<=MEMORY_SIZE was changed to
--		  CONV_INTEGER(low_address)<=MEMORY_SIZE-3
-- 		This avoids an error that freezes the simulation when the
--		   ALU contains a large number (>65533) in its output 
--		   immediately before an LW or SW instruction.
-------------------------------------------------------------------------

library IEEE;
use IEEE.Std_Logic_1164.all;
use std.textio.all;
package aux_functions is  

   subtype wires32  is std_logic_vector(31 downto 0);
   subtype wires16  is std_logic_vector(15 downto 0);
   subtype wires8   is std_logic_vector( 7 downto 0);
   subtype wires4   is std_logic_vector( 3 downto 0);

   -- definição do tipo 'memory', que será utilizado para as memórias de dados/instruções
   constant MEMORY_SIZE : integer := 2048;     
   type memory is array (0 to MEMORY_SIZE) of wires8;

   constant TAM_LINHA : integer := 200;
   
   function CONV_VECTOR( letra : string(1 to TAM_LINHA);  pos: integer ) return std_logic_vector;
	
	procedure readFileLine(file in_file: TEXT; outStrLine: out string);
   
end aux_functions;

package body aux_functions is

  --
  -- converte um caracter de uma dada linha em um std_logic_vector
  --
  function CONV_VECTOR( letra:string(1 to TAM_LINHA);  pos: integer ) return std_logic_vector is         
     variable bin: wires4;
   begin
      case (letra(pos)) is  
              when '0' => bin := "0000";
              when '1' => bin := "0001";
              when '2' => bin := "0010";
              when '3' => bin := "0011";
              when '4' => bin := "0100";
              when '5' => bin := "0101";
              when '6' => bin := "0110";
              when '7' => bin := "0111";
              when '8' => bin := "1000";
              when '9' => bin := "1001";
              when 'A' | 'a' => bin := "1010";
              when 'B' | 'b' => bin := "1011";
              when 'C' | 'c' => bin := "1100";
              when 'D' | 'd' => bin := "1101";
              when 'E' | 'e' => bin := "1110";
              when 'F' | 'f' => bin := "1111";
              when others =>  bin := "0000";  
      end case;
     return bin;
  end CONV_VECTOR;

  procedure readFileLine(file in_file: TEXT; 
					      outStrLine: out string) is
		
		variable localLine: line;
		variable localChar:  character;
		variable isString: 	boolean;
			
	begin
				
		 readline(in_file, localLine);

		 for i in outStrLine'range loop
			 outStrLine(i) := ' ';
		 end loop;   

		 for i in outStrLine'range loop
			read(localLine, localChar, isString);
			outStrLine(i) := localChar;
			if not isString then -- found end of line
				exit;
			end if;   
		 end loop; 
						 
	end readFileLine;
	
end aux_functions;     

--------------------------------------------------------------------------
-- Module implementing a behavioral model of an ASYNCHRONOUS INTERFACE RAM
--------------------------------------------------------------------------
library IEEE;
use ieee.std_logic_1164.all;
use ieee.STD_LOGIC_UNSIGNED.all;
use std.textio.all;
use work.aux_functions.all;

entity RAM_mem is
      generic(  START_ADDRESS: wires32 := (others=>'0')  );
      port( ce_n, we_n, oe_n, bw: in std_logic;    address: in wires32;   data: inout wires32);
end RAM_mem;

architecture RAM_mem of RAM_mem is 
   signal RAM : memory;
   signal tmp_address: wires32;
   alias  low_address: wires16 is tmp_address(15 downto 0);    --  baixa para 16 bits devido ao CONV_INTEGER --
begin     

   tmp_address <= address - START_ADDRESS;   --  offset do endereçamento  -- 
   
   -- writes in memory ASYNCHRONOUSLY  -- LITTLE ENDIAN -------------------
   process(ce_n, we_n, low_address) -- Modification in 16/05/2012 for monocycle processors only,
     begin
       if ce_n='0' and we_n='0' then
          if CONV_INTEGER(low_address)>=0 and CONV_INTEGER(low_address)<=MEMORY_SIZE-3 then
               if bw='1' then
                   RAM(CONV_INTEGER(low_address+3)) <= data(31 downto 24);
                   RAM(CONV_INTEGER(low_address+2)) <= data(23 downto 16);
                   RAM(CONV_INTEGER(low_address+1)) <= data(15 downto  8);
               end if;
               RAM(CONV_INTEGER(low_address  )) <= data( 7 downto  0); 
          end if;
         end if;   
    end process;   
    
   -- read from memory
   process(ce_n, oe_n, low_address)
     begin
       if ce_n='0' and oe_n='0' and
          CONV_INTEGER(low_address)>=0 and CONV_INTEGER(low_address)<=MEMORY_SIZE-3 then
            data(31 downto 24) <= RAM(CONV_INTEGER(low_address+3));
            data(23 downto 16) <= RAM(CONV_INTEGER(low_address+2));
            data(15 downto  8) <= RAM(CONV_INTEGER(low_address+1));
            data( 7 downto  0) <= RAM(CONV_INTEGER(low_address  ));
        else
            data(31 downto 24) <= (others=>'Z');
            data(23 downto 16) <= (others=>'Z');
            data(15 downto  8) <= (others=>'Z');
            data( 7 downto  0) <= (others=>'Z');
        end if;
   end process;   

end RAM_mem;


-------------------------------------------------------------------------
-- pt_br: IMPLEMENTACAO DO MODULO DE PERIFERICO(TB)
-- en_us: IMPLEMENTATION OF THE PERIPHERAL MODULE(TB)
-------------------------------------------------------------------------
library ieee;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;          
use IEEE.std_logic_arith.all;

entity Peripheral is 
port(
      txd : out std_logic;
      rxd : in std_logic;

      clock : in std_logic;
      reset : in std_logic
    );
end entity;

architecture Peripheral of Peripheral is
    signal txd_data: std_logic_vector(9 downto 0);
    
    signal rxd_data1: std_logic_vector(9 downto 0); --start/byte/stop
    signal rxd_data2: std_logic_vector(9 downto 0); --start/byte/stop
    -- pt_br: Estados da FSM 
    -- en_us: FSM States
    type State is (A,B,C,D,E);
    -- pt_br: estado atual
    -- en_us: current state
    signal st : State;

    -- pt_br: nao esta sendo utilizada, o intervalo de tempo e colocado pelo sistema
    -- en_us: it isn't beeing used, the time interval is beeing generated by the system
    --constant bps : time := 8.68 us; -- 115.200 bps

    signal txd_count: std_logic_vector(8 downto 0) := (others => '0');

    -- pt_br: Sinais de depuracao
    -- en_us: Debugging signal

    --signal debug: std_logic := '0';
    --signal debug2: std_logic := '0';
    --signal debug3: std_logic := '0';

begin
  
Peripheral_FSM:  process(clock,reset)
  begin
    if reset = '1' then
      rxd_data1 <= (others => '1');
      rxd_data2 <= (others => '1');
      txd_data <= (others => '1');
    elsif clock = '1' and clock'event then
      case st is
          -- pt_br: 0x55 configura MEF de autobaud
          -- en_us: 0x55 configure MEF autobaud
          when A =>
            txd_data <= '1' & "01010101" & '0';
            txd_count <= (8 => '0', others => '1');
            st <= E;

          -- pt_br: espera receber o primeiro dado
          -- en_us: wait to receive first data
          when B =>
            --debug <= '1';
            -- pt_br: ele verifica em 1, pois leva 1 ciclo p/ receber o ultimo valor
            -- en_us: it verifies (1) because it takes 1 cycle to receive the last value
            if rxd_data1(1) = '0' then
              st <= C;
            end if;
            rxd_data1 <= rxd & rxd_data1(9 downto 1);
          -- pt_br: espera receber o segundo dado
          -- en_us: wait to receive second data
          when C =>
            --debug3 <= '1';

            -- pt_br: para
            -- en_us: stop
            if rxd_data2(0) = '0' then
              st <= D;
            else
              rxd_data2 <= rxd & rxd_data2(9 downto 1);  
            end if;
          -- pt_br: soma os valores e manda o bit '0' p/ iniciar
          -- en_us: sum two values and send 0 bit to start
          when D => 
            txd_data <= '1' & rxd_data1(8 downto 1) + rxd_data2(8 downto 1) & '0';
            txd_count <= (8 => '0', others => '1');
            st <= E;
          -- pt_br: manda os outros 9 bits (dado e '1' p/ terminar)
          -- en_us: send the other 9 bits (data and '1' to end)
          when E => 
            txd_data <= '1' & txd_data(9 downto 1);
            txd_count <= '0' & txd_count(8 downto 1);
            -- pt_br: acabou !
            -- en_us: it's over !
            if txd_count(0) = '0' then
              -- pt_br: zera os 2
              -- en_us: clear both registers
              rxd_data1 <= (others => '1');
              rxd_data2 <= (others => '1');
              st <= B;
            end if;
      end case;
    end if;
  end process;

-- pt_br: O txd sendo enviado, txd_data eh atualizada em rising edge
-- en_us: txd beeing sent, txd_data is updated in rising edge
txd <= txd_data(0);

end Peripheral;
-------------------------------------------------------------------------
-- pt_br: IMPLEMENTACAO DO TESTBENCH DO SISTEMA
-- en_us: IMPLEMENTATION OF THE SYSTEM TESTBENCH 
-------------------------------------------------------------------------
library ieee;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;          
use STD.TEXTIO.all;
use work.aux_functions.all;
entity system_tb is
end system_tb;

architecture system_tb of system_tb is
  ----------------------------------------------------
  ------ pt_br: Sinais do Periferico
  ------ en_us: Peripheral Signals
  ----------------------------------------------------
  signal Pclock,Preset : std_logic;
  ----------------------------------------------------
  ------ pt_br: Sinais da Interface Serial C/ Peripheral
  ------ en_us: Signas of the Serial Interface W/ Peripheral
  ----------------------------------------------------
  signal rxd,txd : std_logic;
  ----------------------------------------------------
  ------ pt_br: Sinais da Logica de Cola C/ Interface Serial
  ------ en_us: Glue logic signal W/ Serial Interface
  ----------------------------------------------------

  signal rx_data : wires8 := (others => '0');
  signal rx_start, rx_busy : std_logic;

  signal tx_data : wires8 := (others => '0');
  signal tx_av : std_logic;
  ----------------------------------------------------
  ------ pt_br: Sinal da Logica de Cola C/ Memoria(TB) e CPU(HW)
  ------ en_us: Glue Logic signals W/ Memory(TB) and CPU(HW)
  ----------------------------------------------------
  signal GLaddress : wires32 := (others => '0');
  signal GLdata : wires32 := (others => '0');

  ----------------------------------------------------
  ------ pt_br: Sinais da CPU
  ------ en_us: CPU Signals
  ----------------------------------------------------
  signal Dadress, Ddata, Iadress, Idata,
         i_cpu_address, d_cpu_address, data_cpu,
         tb_add, tb_data : wires32 := (others => '0' );
  
  signal Dce_n, Dwe_n, Doe_n, Ice_n, Iwe_n, Ioe_n, ck, rst, rstCPU,
         go_i, go_d, ce, rw, bw: std_logic;
  
  -----------------------------------------------------------------

  -- pt_br: Arquivo gerado pelo simulador MARS que sera utilizado 
  -- para carregar as instrucoes e memoria de dados. Dependendo do
  -- sistema em que tal simulacao ocorre talvez seja necessario 
  -- adicionar todo o caminho ate o arquivo.

  -- en_us: File generated by MARS Simulator which will be used to
  -- load the instructions and data memory. Depending on the system
  -- on which the simulation will occur, it may be necessary to
  -- write the full path to the file.
  file ARQ : TEXT open READ_MODE is "softwareText.txt";
  
  -----------------------------------------------------------------

begin 
  -------------------------------------------------
    -- pt_br: Memoria de Dados
    -- en_us: Data Memory
  Data_mem: entity work.RAM_mem 
    generic map( START_ADDRESS => x"10010000" )
    port map(
      ce_n => Dce_n,
      we_n => Dwe_n,
      oe_n => Doe_n,
      bw => bw,
      address => Dadress,
      data => Ddata
    );
    -- pt_br: Memoria de Instrucoes
    -- en_us: Instruction Memory
  Instr_mem: entity work.RAM_mem 
    generic map( START_ADDRESS => x"00400000" )
    port map(
      ce_n =>Ice_n,
      we_n =>Iwe_n,
      oe_n =>Ioe_n,
      bw => '1',
      address => Iadress,
      data => Idata
    );

  -------------------------------------------------
  -- pt_br: Logica de Cola
  -- en_us: Glue Logic
  glueLogic: entity work.glueLogic
    port map(
      clock => ck,
      reset => rstCPU,
      tx_data => tx_data,
      tx_av => tx_av,
      rx_data => rx_data,
      rx_start => rx_start,
      rx_busy => rx_busy,
      data => GLdata,
      ce => ce,
      rw => rw,
      address => GLaddress
    );  
  --------------------------------------------------
  -- pt_br: Interface Serial
  -- en_us: Serial Interface
  serialInterface: entity work.serialinterface
    port map(
        clock => ck,
        reset => rstCPU,
        rxd => rxd,
        txd => txd,
        rx_data => rx_data,
        rx_start => rx_start,
        rx_busy => rx_busy,
        tx_data => tx_data,
        tx_av => tx_av
    );

    -- pt_br: Periferico
    -- en_us: Peripheral
    peripheral: entity work.Peripheral
    port map(
        txd => txd,
        rxd => rxd,
        clock => Pclock,
        reset => Preset
    );

  -------------------------------------
    -- pt_br: O proprio processador
    -- en_us: The CPU itself
    cpu: entity work.MIPS_MCS
      port map(
        clock => ck,
        reset => rstCPU,
        i_address => i_cpu_address,
        instruction => Idata,
        ce => ce,
        rw => rw,
        bw => bw,
        d_address => d_cpu_address,
        data => data_cpu
      );


    -- data memory signals --------------------------------------------------------
    Dce_n <= '0' when (ce='1' and rstCPU/='1') or go_d='1' else '1'; -- Bug corrected here in 16/05/2012
    
    Doe_n <= '0' when (ce='1' and rw='1')             else '1';       
    Dwe_n <= '0' when (ce='1' and rw='0') or go_d='1' else '1';    

    Dadress <= tb_add  when rstCPU='1' else d_cpu_address;
    
    Ddata   <= tb_data when rstCPU='1' else data_cpu when (ce='1' and rw='0') else (others=>'Z'); 
    
    -- pt_br: Recebe da Logica de Cola quando o endereco for um dos 10008...
    -- Recebe da memoria de dados caso seja um endereco dela 1001...

    -- en_us: Receives from the Glue Logic when the adress matches 10008...
    -- Receives from the data memory if the address matches 1001...
    data_cpu <= Ddata when (ce = '1' and rw = '1') and d_cpu_address(31 downto 16) = x"1001" else
                GLdata when (ce = '1' and rw = '1') and d_cpu_address(31 downto 12) = x"10008"
                else (others => 'Z');

    
    -- instructions memory signals --------------------------------------------------------
    Ice_n <= '0';                               
    -- pt_br: impede leitura enquanto está escrevendo                               
    -- en_us: block reading while its writign
    Ioe_n <= '1' when rstCPU='1' else '0';   
    -- pt_br: impede escrita durante a leitura do arquivo    
    -- en_us: blocks write while the file is beeing read
    Iwe_n <= '0' when go_i='1'   else '1';   
    
    Iadress <= tb_add  when rstCPU='1' else i_cpu_address;
    Idata   <= tb_data when rstCPU='1' else (others => 'Z'); 

    -- pt_br: Endereco da Logica de Cola
    -- en_us: Glue Logic Address
    GLaddress <= d_cpu_address when rstCPU = '0' else (others => 'Z');

    
    -- pt_br: Dado da logica de cola
    -- en_us: Glue Logic Data
    GLdata <= data_cpu when rstCPU = '0' else (others => 'Z');
    

    -- pt_br: Gera o Clock do periferico --
    -- en_us: Generates Peripheral Clock
    process
      begin
        Pclock <= '1', '0' after 4.34 us;
        wait for 8.68 us;
    end process;

    Preset <= '1', '0' after 8.68 us;


--------------------------------------------------------------------------------------------

  rst <='1', '0' after 15 ns;       -- generates the reset signal 


  process                          -- generates the clock signal 
      begin
      ck <= '1', '0' after 10 ns;
      wait for 20 ns;
  end process;

    ----------------------------------------------------------------------------
    -- this process loads the instruction memory and the data memory during reset
    --
    --
    --   O PROCESSO ABAIXO EH UMA PARSER PARA LER CODIGO GERADO PELO SPIM NO
    --   SEGUINTE FORMATO:
    --
    --      Text Segment
    --      [0x00400000]        0x3c011001  lui $1, 4097 [d2]               ; 16: la    $t0, d2
    --      [0x00400004]        0x34280004  ori $8, $1, 4 [d2]
    --      [0x00400008]        0x8d080000  lw $8, 0($8)                    ; 17: lw    $t0,0($t0)
    --      .....
    --      [0x00400048]        0x0810000f  j 0x0040003c [loop]             ; 30: j     loop
    --      [0x0040004c]        0x01284821  addu $9, $9, $8                 ; 32: addu $t1, $t1, $t0
    --      [0x00400050]        0x08100014  j 0x00400050 [x]                ; 34: j     x
    --      Data Segment
    --      [0x10010000]                        0x0000faaa  0x00000083  0x00000000  0x00000000
    --
    ----------------------------------------------------------------------------
    process
        variable ARQ_LINE : LINE;
        variable line_arq : string(1 to TAM_LINHA);
        variable code     : boolean;
        variable i, address_flag : integer;
    begin  
        go_i <= '0';
        go_d <= '0';
        rstCPU <= '1';           -- hold the processor during file reading
        code:=true;              -- default value of code is 1 (CODE)
                                 
        wait until rst = '1';
        
        while NOT (endfile(ARQ)) loop    -- INICIO DA LEITURA DO ARQUIVO CONTENDO INSTRUCAO E DADOS -----
            --readline(ARQ, ARQ_LINE);      
            --read(ARQ_LINE, line_arq(1 to  ARQ_LINE'length) );
        readFileLine(ARQ, line_arq);
                        
            if line_arq(1 to 12)="Text Segment" then 
                   code:=true;                     -- code 
            elsif line_arq(1 to 12)="Data Segment" then
                   code:=false;                    -- data 
            else 
               i := 1;                                  -- LEITORA DE LINHA - analizar o loop abaixo para compreender 
               address_flag := 0;                       -- para INSTRUCAO é um para (end,inst)
                                                        -- para DADO aceita (end, dado 0, dado 1, dado 2 ....)
               loop                                     
                  if line_arq(i) = '0' and line_arq(i+1) = 'x' then      -- encontrou indicacao de numero hexa: '0x'
                         i := i + 2;
                         if address_flag=0 then
                               for w in 0 to 7 loop
                                   tb_add( (31-w*4) downto (32-(w+1)*4))  <= CONV_VECTOR(line_arq,i+w);
                               end loop;    
                               i := i + 8; 
                               address_flag := 1;
                         else
                               for w in 0 to 7 loop
                                   tb_data( (31-w*4) downto (32-(w+1)*4))  <= CONV_VECTOR(line_arq,i+w);
                               end loop;    
                               i := i + 8;
                               
                               wait for 0.1 ns;
                               
                               if code=true then go_i <= '1';    -- the go_i signal enables instruction memory writing
                                            else go_d <= '1';    -- the go_d signal enables data memory writing
                               end if; 
                               
                               wait for 0.1 ns;
                               
                               tb_add <= tb_add + 4;       -- *great!* consigo ler mais de uma word por linha!
                               go_i <= '0';
                               go_d <= '0'; 
                               
                               address_flag := 2;    -- sinaliza que ja leu o conteudo do endereco;

                         end if;
                  end if;
                  i := i + 1;
                  
                  -- sai da linha quando chegou no seu final OU ja leu par(endereço, instrucao) no caso de codigo
                  exit when i=TAM_LINHA or (code=true and address_flag=2);
               end loop;
            end if;
            
        end loop;                        -- FINAL DA LEITURA DO ARQUIVO CONTENDO INSTRUCAO E DADOS -----
        
        rstCPU <= '0' after 2 ns;   -- release the processor to execute
        wait for 4 ns;   -- To activate the RST CPU signal
        wait until rst = '1';  -- to Hold again!
        
    end process;

end system_tb;